/*************************************************************

    Filename    : simple_soc_test_lib.sv
    Author      : yyl
    Description : 
    Creat Time  : 2025-03-15 02:21:49
    Modify Time : 2025-03-15 02:21:49

*************************************************************/
`ifndef SIMPLE_SOC_TEST_LIB__SV
`define SIMPLE_SOC_TEST_LIB__SV

`soc_create_test(debug,0)

`endif
